module fixed_mult
#(
  parameter L = 16
)
(
  input wire [L - 1: 0] a,
  input wire [L - 1: 0] b,
  output wire [L - 1: 0] c
);

endmodule
