`timescale 1ns/1ps

module fixed_mult_tb();

endmodule
